/*==========================================================*/

//generate year month day signals output to display moudle

/*==========================================================*/
module example (
    input clk,    // Clock
    input clk_en, // Clock Enable
    input rst_n,  // Asynchronous reset active low
    
);





/***********************************************************/
endmodule
/*==========================================================*/
